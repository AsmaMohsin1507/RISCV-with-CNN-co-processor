magic
tech gf180mcuC
magscale 1 5
timestamp 1670049064
<< obsm1 >>
rect 672 855 59304 58561
<< metal2 >>
rect 336 59600 392 59900
rect 1008 59600 1064 59900
rect 1680 59600 1736 59900
rect 2016 59600 2072 59900
rect 2688 59600 2744 59900
rect 3360 59600 3416 59900
rect 4032 59600 4088 59900
rect 4368 59600 4424 59900
rect 5040 59600 5096 59900
rect 5712 59600 5768 59900
rect 6048 59600 6104 59900
rect 6720 59600 6776 59900
rect 7392 59600 7448 59900
rect 8064 59600 8120 59900
rect 8400 59600 8456 59900
rect 9072 59600 9128 59900
rect 9744 59600 9800 59900
rect 10080 59600 10136 59900
rect 10752 59600 10808 59900
rect 11424 59600 11480 59900
rect 12096 59600 12152 59900
rect 12432 59600 12488 59900
rect 13104 59600 13160 59900
rect 13776 59600 13832 59900
rect 14448 59600 14504 59900
rect 14784 59600 14840 59900
rect 15456 59600 15512 59900
rect 16128 59600 16184 59900
rect 16464 59600 16520 59900
rect 17136 59600 17192 59900
rect 17808 59600 17864 59900
rect 18480 59600 18536 59900
rect 18816 59600 18872 59900
rect 19488 59600 19544 59900
rect 20160 59600 20216 59900
rect 20496 59600 20552 59900
rect 21168 59600 21224 59900
rect 21840 59600 21896 59900
rect 22512 59600 22568 59900
rect 22848 59600 22904 59900
rect 23520 59600 23576 59900
rect 24192 59600 24248 59900
rect 24864 59600 24920 59900
rect 25200 59600 25256 59900
rect 25872 59600 25928 59900
rect 26544 59600 26600 59900
rect 26880 59600 26936 59900
rect 27552 59600 27608 59900
rect 28224 59600 28280 59900
rect 28896 59600 28952 59900
rect 29232 59600 29288 59900
rect 29904 59600 29960 59900
rect 30576 59600 30632 59900
rect 30912 59600 30968 59900
rect 31584 59600 31640 59900
rect 32256 59600 32312 59900
rect 32928 59600 32984 59900
rect 33264 59600 33320 59900
rect 33936 59600 33992 59900
rect 34608 59600 34664 59900
rect 34944 59600 35000 59900
rect 35616 59600 35672 59900
rect 36288 59600 36344 59900
rect 36960 59600 37016 59900
rect 37296 59600 37352 59900
rect 37968 59600 38024 59900
rect 38640 59600 38696 59900
rect 39312 59600 39368 59900
rect 39648 59600 39704 59900
rect 40320 59600 40376 59900
rect 40992 59600 41048 59900
rect 41328 59600 41384 59900
rect 42000 59600 42056 59900
rect 42672 59600 42728 59900
rect 43344 59600 43400 59900
rect 43680 59600 43736 59900
rect 44352 59600 44408 59900
rect 45024 59600 45080 59900
rect 45360 59600 45416 59900
rect 46032 59600 46088 59900
rect 46704 59600 46760 59900
rect 47376 59600 47432 59900
rect 47712 59600 47768 59900
rect 48384 59600 48440 59900
rect 49056 59600 49112 59900
rect 49728 59600 49784 59900
rect 50064 59600 50120 59900
rect 50736 59600 50792 59900
rect 51408 59600 51464 59900
rect 51744 59600 51800 59900
rect 52416 59600 52472 59900
rect 53088 59600 53144 59900
rect 53760 59600 53816 59900
rect 54096 59600 54152 59900
rect 54768 59600 54824 59900
rect 55440 59600 55496 59900
rect 55776 59600 55832 59900
rect 56448 59600 56504 59900
rect 57120 59600 57176 59900
rect 57792 59600 57848 59900
rect 58128 59600 58184 59900
rect 58800 59600 58856 59900
rect 59472 59600 59528 59900
rect 59808 59600 59864 59900
rect 0 100 56 400
rect 336 100 392 400
rect 1008 100 1064 400
rect 1680 100 1736 400
rect 2016 100 2072 400
rect 2688 100 2744 400
rect 3360 100 3416 400
rect 4032 100 4088 400
rect 4368 100 4424 400
rect 5040 100 5096 400
rect 5712 100 5768 400
rect 6048 100 6104 400
rect 6720 100 6776 400
rect 7392 100 7448 400
rect 8064 100 8120 400
rect 8400 100 8456 400
rect 9072 100 9128 400
rect 9744 100 9800 400
rect 10080 100 10136 400
rect 10752 100 10808 400
rect 11424 100 11480 400
rect 12096 100 12152 400
rect 12432 100 12488 400
rect 13104 100 13160 400
rect 13776 100 13832 400
rect 14448 100 14504 400
rect 14784 100 14840 400
rect 15456 100 15512 400
rect 16128 100 16184 400
rect 16464 100 16520 400
rect 17136 100 17192 400
rect 17808 100 17864 400
rect 18480 100 18536 400
rect 18816 100 18872 400
rect 19488 100 19544 400
rect 20160 100 20216 400
rect 20496 100 20552 400
rect 21168 100 21224 400
rect 21840 100 21896 400
rect 22512 100 22568 400
rect 22848 100 22904 400
rect 23520 100 23576 400
rect 24192 100 24248 400
rect 24864 100 24920 400
rect 25200 100 25256 400
rect 25872 100 25928 400
rect 26544 100 26600 400
rect 26880 100 26936 400
rect 27552 100 27608 400
rect 28224 100 28280 400
rect 28896 100 28952 400
rect 29232 100 29288 400
rect 29904 100 29960 400
rect 30576 100 30632 400
rect 30912 100 30968 400
rect 31584 100 31640 400
rect 32256 100 32312 400
rect 32928 100 32984 400
rect 33264 100 33320 400
rect 33936 100 33992 400
rect 34608 100 34664 400
rect 34944 100 35000 400
rect 35616 100 35672 400
rect 36288 100 36344 400
rect 36960 100 37016 400
rect 37296 100 37352 400
rect 37968 100 38024 400
rect 38640 100 38696 400
rect 39312 100 39368 400
rect 39648 100 39704 400
rect 40320 100 40376 400
rect 40992 100 41048 400
rect 41328 100 41384 400
rect 42000 100 42056 400
rect 42672 100 42728 400
rect 43344 100 43400 400
rect 43680 100 43736 400
rect 44352 100 44408 400
rect 45024 100 45080 400
rect 45360 100 45416 400
rect 46032 100 46088 400
rect 46704 100 46760 400
rect 47376 100 47432 400
rect 47712 100 47768 400
rect 48384 100 48440 400
rect 49056 100 49112 400
rect 49728 100 49784 400
rect 50064 100 50120 400
rect 50736 100 50792 400
rect 51408 100 51464 400
rect 51744 100 51800 400
rect 52416 100 52472 400
rect 53088 100 53144 400
rect 53760 100 53816 400
rect 54096 100 54152 400
rect 54768 100 54824 400
rect 55440 100 55496 400
rect 55776 100 55832 400
rect 56448 100 56504 400
rect 57120 100 57176 400
rect 57792 100 57848 400
rect 58128 100 58184 400
rect 58800 100 58856 400
rect 59472 100 59528 400
<< obsm2 >>
rect 14 59570 306 59911
rect 422 59570 978 59911
rect 1094 59570 1650 59911
rect 1766 59570 1986 59911
rect 2102 59570 2658 59911
rect 2774 59570 3330 59911
rect 3446 59570 4002 59911
rect 4118 59570 4338 59911
rect 4454 59570 5010 59911
rect 5126 59570 5682 59911
rect 5798 59570 6018 59911
rect 6134 59570 6690 59911
rect 6806 59570 7362 59911
rect 7478 59570 8034 59911
rect 8150 59570 8370 59911
rect 8486 59570 9042 59911
rect 9158 59570 9714 59911
rect 9830 59570 10050 59911
rect 10166 59570 10722 59911
rect 10838 59570 11394 59911
rect 11510 59570 12066 59911
rect 12182 59570 12402 59911
rect 12518 59570 13074 59911
rect 13190 59570 13746 59911
rect 13862 59570 14418 59911
rect 14534 59570 14754 59911
rect 14870 59570 15426 59911
rect 15542 59570 16098 59911
rect 16214 59570 16434 59911
rect 16550 59570 17106 59911
rect 17222 59570 17778 59911
rect 17894 59570 18450 59911
rect 18566 59570 18786 59911
rect 18902 59570 19458 59911
rect 19574 59570 20130 59911
rect 20246 59570 20466 59911
rect 20582 59570 21138 59911
rect 21254 59570 21810 59911
rect 21926 59570 22482 59911
rect 22598 59570 22818 59911
rect 22934 59570 23490 59911
rect 23606 59570 24162 59911
rect 24278 59570 24834 59911
rect 24950 59570 25170 59911
rect 25286 59570 25842 59911
rect 25958 59570 26514 59911
rect 26630 59570 26850 59911
rect 26966 59570 27522 59911
rect 27638 59570 28194 59911
rect 28310 59570 28866 59911
rect 28982 59570 29202 59911
rect 29318 59570 29874 59911
rect 29990 59570 30546 59911
rect 30662 59570 30882 59911
rect 30998 59570 31554 59911
rect 31670 59570 32226 59911
rect 32342 59570 32898 59911
rect 33014 59570 33234 59911
rect 33350 59570 33906 59911
rect 34022 59570 34578 59911
rect 34694 59570 34914 59911
rect 35030 59570 35586 59911
rect 35702 59570 36258 59911
rect 36374 59570 36930 59911
rect 37046 59570 37266 59911
rect 37382 59570 37938 59911
rect 38054 59570 38610 59911
rect 38726 59570 39282 59911
rect 39398 59570 39618 59911
rect 39734 59570 40290 59911
rect 40406 59570 40962 59911
rect 41078 59570 41298 59911
rect 41414 59570 41970 59911
rect 42086 59570 42642 59911
rect 42758 59570 43314 59911
rect 43430 59570 43650 59911
rect 43766 59570 44322 59911
rect 44438 59570 44994 59911
rect 45110 59570 45330 59911
rect 45446 59570 46002 59911
rect 46118 59570 46674 59911
rect 46790 59570 47346 59911
rect 47462 59570 47682 59911
rect 47798 59570 48354 59911
rect 48470 59570 49026 59911
rect 49142 59570 49698 59911
rect 49814 59570 50034 59911
rect 50150 59570 50706 59911
rect 50822 59570 51378 59911
rect 51494 59570 51714 59911
rect 51830 59570 52386 59911
rect 52502 59570 53058 59911
rect 53174 59570 53730 59911
rect 53846 59570 54066 59911
rect 54182 59570 54738 59911
rect 54854 59570 55410 59911
rect 55526 59570 55746 59911
rect 55862 59570 56418 59911
rect 56534 59570 57090 59911
rect 57206 59570 57762 59911
rect 57878 59570 58098 59911
rect 58214 59570 58770 59911
rect 58886 59570 59442 59911
rect 59558 59570 59626 59911
rect 14 430 59626 59570
rect 86 400 306 430
rect 422 400 978 430
rect 1094 400 1650 430
rect 1766 400 1986 430
rect 2102 400 2658 430
rect 2774 400 3330 430
rect 3446 400 4002 430
rect 4118 400 4338 430
rect 4454 400 5010 430
rect 5126 400 5682 430
rect 5798 400 6018 430
rect 6134 400 6690 430
rect 6806 400 7362 430
rect 7478 400 8034 430
rect 8150 400 8370 430
rect 8486 400 9042 430
rect 9158 400 9714 430
rect 9830 400 10050 430
rect 10166 400 10722 430
rect 10838 400 11394 430
rect 11510 400 12066 430
rect 12182 400 12402 430
rect 12518 400 13074 430
rect 13190 400 13746 430
rect 13862 400 14418 430
rect 14534 400 14754 430
rect 14870 400 15426 430
rect 15542 400 16098 430
rect 16214 400 16434 430
rect 16550 400 17106 430
rect 17222 400 17778 430
rect 17894 400 18450 430
rect 18566 400 18786 430
rect 18902 400 19458 430
rect 19574 400 20130 430
rect 20246 400 20466 430
rect 20582 400 21138 430
rect 21254 400 21810 430
rect 21926 400 22482 430
rect 22598 400 22818 430
rect 22934 400 23490 430
rect 23606 400 24162 430
rect 24278 400 24834 430
rect 24950 400 25170 430
rect 25286 400 25842 430
rect 25958 400 26514 430
rect 26630 400 26850 430
rect 26966 400 27522 430
rect 27638 400 28194 430
rect 28310 400 28866 430
rect 28982 400 29202 430
rect 29318 400 29874 430
rect 29990 400 30546 430
rect 30662 400 30882 430
rect 30998 400 31554 430
rect 31670 400 32226 430
rect 32342 400 32898 430
rect 33014 400 33234 430
rect 33350 400 33906 430
rect 34022 400 34578 430
rect 34694 400 34914 430
rect 35030 400 35586 430
rect 35702 400 36258 430
rect 36374 400 36930 430
rect 37046 400 37266 430
rect 37382 400 37938 430
rect 38054 400 38610 430
rect 38726 400 39282 430
rect 39398 400 39618 430
rect 39734 400 40290 430
rect 40406 400 40962 430
rect 41078 400 41298 430
rect 41414 400 41970 430
rect 42086 400 42642 430
rect 42758 400 43314 430
rect 43430 400 43650 430
rect 43766 400 44322 430
rect 44438 400 44994 430
rect 45110 400 45330 430
rect 45446 400 46002 430
rect 46118 400 46674 430
rect 46790 400 47346 430
rect 47462 400 47682 430
rect 47798 400 48354 430
rect 48470 400 49026 430
rect 49142 400 49698 430
rect 49814 400 50034 430
rect 50150 400 50706 430
rect 50822 400 51378 430
rect 51494 400 51714 430
rect 51830 400 52386 430
rect 52502 400 53058 430
rect 53174 400 53730 430
rect 53846 400 54066 430
rect 54182 400 54738 430
rect 54854 400 55410 430
rect 55526 400 55746 430
rect 55862 400 56418 430
rect 56534 400 57090 430
rect 57206 400 57762 430
rect 57878 400 58098 430
rect 58214 400 58770 430
rect 58886 400 59442 430
rect 59558 400 59626 430
<< metal3 >>
rect 100 59808 400 59864
rect 100 59472 400 59528
rect 59600 59472 59900 59528
rect 100 58800 400 58856
rect 59600 58800 59900 58856
rect 100 58128 400 58184
rect 59600 58128 59900 58184
rect 100 57792 400 57848
rect 59600 57792 59900 57848
rect 100 57120 400 57176
rect 59600 57120 59900 57176
rect 100 56448 400 56504
rect 59600 56448 59900 56504
rect 100 55776 400 55832
rect 59600 55776 59900 55832
rect 100 55440 400 55496
rect 59600 55440 59900 55496
rect 100 54768 400 54824
rect 59600 54768 59900 54824
rect 100 54096 400 54152
rect 59600 54096 59900 54152
rect 100 53760 400 53816
rect 59600 53760 59900 53816
rect 100 53088 400 53144
rect 59600 53088 59900 53144
rect 100 52416 400 52472
rect 59600 52416 59900 52472
rect 100 51744 400 51800
rect 59600 51744 59900 51800
rect 100 51408 400 51464
rect 59600 51408 59900 51464
rect 100 50736 400 50792
rect 59600 50736 59900 50792
rect 100 50064 400 50120
rect 59600 50064 59900 50120
rect 100 49728 400 49784
rect 59600 49728 59900 49784
rect 100 49056 400 49112
rect 59600 49056 59900 49112
rect 100 48384 400 48440
rect 59600 48384 59900 48440
rect 100 47712 400 47768
rect 59600 47712 59900 47768
rect 100 47376 400 47432
rect 59600 47376 59900 47432
rect 100 46704 400 46760
rect 59600 46704 59900 46760
rect 100 46032 400 46088
rect 59600 46032 59900 46088
rect 100 45360 400 45416
rect 59600 45360 59900 45416
rect 100 45024 400 45080
rect 59600 45024 59900 45080
rect 100 44352 400 44408
rect 59600 44352 59900 44408
rect 100 43680 400 43736
rect 59600 43680 59900 43736
rect 100 43344 400 43400
rect 59600 43344 59900 43400
rect 100 42672 400 42728
rect 59600 42672 59900 42728
rect 100 42000 400 42056
rect 59600 42000 59900 42056
rect 100 41328 400 41384
rect 59600 41328 59900 41384
rect 100 40992 400 41048
rect 59600 40992 59900 41048
rect 100 40320 400 40376
rect 59600 40320 59900 40376
rect 100 39648 400 39704
rect 59600 39648 59900 39704
rect 100 39312 400 39368
rect 59600 39312 59900 39368
rect 100 38640 400 38696
rect 59600 38640 59900 38696
rect 100 37968 400 38024
rect 59600 37968 59900 38024
rect 100 37296 400 37352
rect 59600 37296 59900 37352
rect 100 36960 400 37016
rect 59600 36960 59900 37016
rect 100 36288 400 36344
rect 59600 36288 59900 36344
rect 100 35616 400 35672
rect 59600 35616 59900 35672
rect 100 34944 400 35000
rect 59600 34944 59900 35000
rect 100 34608 400 34664
rect 59600 34608 59900 34664
rect 100 33936 400 33992
rect 59600 33936 59900 33992
rect 100 33264 400 33320
rect 59600 33264 59900 33320
rect 100 32928 400 32984
rect 59600 32928 59900 32984
rect 100 32256 400 32312
rect 59600 32256 59900 32312
rect 100 31584 400 31640
rect 59600 31584 59900 31640
rect 100 30912 400 30968
rect 59600 30912 59900 30968
rect 100 30576 400 30632
rect 59600 30576 59900 30632
rect 100 29904 400 29960
rect 59600 29904 59900 29960
rect 100 29232 400 29288
rect 59600 29232 59900 29288
rect 100 28896 400 28952
rect 59600 28896 59900 28952
rect 100 28224 400 28280
rect 59600 28224 59900 28280
rect 100 27552 400 27608
rect 59600 27552 59900 27608
rect 100 26880 400 26936
rect 59600 26880 59900 26936
rect 100 26544 400 26600
rect 59600 26544 59900 26600
rect 100 25872 400 25928
rect 59600 25872 59900 25928
rect 100 25200 400 25256
rect 59600 25200 59900 25256
rect 100 24864 400 24920
rect 59600 24864 59900 24920
rect 100 24192 400 24248
rect 59600 24192 59900 24248
rect 100 23520 400 23576
rect 59600 23520 59900 23576
rect 100 22848 400 22904
rect 59600 22848 59900 22904
rect 100 22512 400 22568
rect 59600 22512 59900 22568
rect 100 21840 400 21896
rect 59600 21840 59900 21896
rect 100 21168 400 21224
rect 59600 21168 59900 21224
rect 100 20496 400 20552
rect 59600 20496 59900 20552
rect 100 20160 400 20216
rect 59600 20160 59900 20216
rect 100 19488 400 19544
rect 59600 19488 59900 19544
rect 100 18816 400 18872
rect 59600 18816 59900 18872
rect 100 18480 400 18536
rect 59600 18480 59900 18536
rect 100 17808 400 17864
rect 59600 17808 59900 17864
rect 100 17136 400 17192
rect 59600 17136 59900 17192
rect 100 16464 400 16520
rect 59600 16464 59900 16520
rect 100 16128 400 16184
rect 59600 16128 59900 16184
rect 100 15456 400 15512
rect 59600 15456 59900 15512
rect 100 14784 400 14840
rect 59600 14784 59900 14840
rect 100 14448 400 14504
rect 59600 14448 59900 14504
rect 100 13776 400 13832
rect 59600 13776 59900 13832
rect 100 13104 400 13160
rect 59600 13104 59900 13160
rect 100 12432 400 12488
rect 59600 12432 59900 12488
rect 100 12096 400 12152
rect 59600 12096 59900 12152
rect 100 11424 400 11480
rect 59600 11424 59900 11480
rect 100 10752 400 10808
rect 59600 10752 59900 10808
rect 100 10080 400 10136
rect 59600 10080 59900 10136
rect 100 9744 400 9800
rect 59600 9744 59900 9800
rect 100 9072 400 9128
rect 59600 9072 59900 9128
rect 100 8400 400 8456
rect 59600 8400 59900 8456
rect 100 8064 400 8120
rect 59600 8064 59900 8120
rect 100 7392 400 7448
rect 59600 7392 59900 7448
rect 100 6720 400 6776
rect 59600 6720 59900 6776
rect 100 6048 400 6104
rect 59600 6048 59900 6104
rect 100 5712 400 5768
rect 59600 5712 59900 5768
rect 100 5040 400 5096
rect 59600 5040 59900 5096
rect 100 4368 400 4424
rect 59600 4368 59900 4424
rect 100 4032 400 4088
rect 59600 4032 59900 4088
rect 100 3360 400 3416
rect 59600 3360 59900 3416
rect 100 2688 400 2744
rect 59600 2688 59900 2744
rect 100 2016 400 2072
rect 59600 2016 59900 2072
rect 100 1680 400 1736
rect 59600 1680 59900 1736
rect 100 1008 400 1064
rect 59600 1008 59900 1064
rect 100 336 400 392
rect 59600 336 59900 392
rect 59600 0 59900 56
<< obsm3 >>
rect 9 59894 59631 59906
rect 9 59778 70 59894
rect 430 59778 59631 59894
rect 9 59558 59631 59778
rect 9 59442 70 59558
rect 430 59442 59570 59558
rect 9 58886 59631 59442
rect 9 58770 70 58886
rect 430 58770 59570 58886
rect 9 58214 59631 58770
rect 9 58098 70 58214
rect 430 58098 59570 58214
rect 9 57878 59631 58098
rect 9 57762 70 57878
rect 430 57762 59570 57878
rect 9 57206 59631 57762
rect 9 57090 70 57206
rect 430 57090 59570 57206
rect 9 56534 59631 57090
rect 9 56418 70 56534
rect 430 56418 59570 56534
rect 9 55862 59631 56418
rect 9 55746 70 55862
rect 430 55746 59570 55862
rect 9 55526 59631 55746
rect 9 55410 70 55526
rect 430 55410 59570 55526
rect 9 54854 59631 55410
rect 9 54738 70 54854
rect 430 54738 59570 54854
rect 9 54182 59631 54738
rect 9 54066 70 54182
rect 430 54066 59570 54182
rect 9 53846 59631 54066
rect 9 53730 70 53846
rect 430 53730 59570 53846
rect 9 53174 59631 53730
rect 9 53058 70 53174
rect 430 53058 59570 53174
rect 9 52502 59631 53058
rect 9 52386 70 52502
rect 430 52386 59570 52502
rect 9 51830 59631 52386
rect 9 51714 70 51830
rect 430 51714 59570 51830
rect 9 51494 59631 51714
rect 9 51378 70 51494
rect 430 51378 59570 51494
rect 9 50822 59631 51378
rect 9 50706 70 50822
rect 430 50706 59570 50822
rect 9 50150 59631 50706
rect 9 50034 70 50150
rect 430 50034 59570 50150
rect 9 49814 59631 50034
rect 9 49698 70 49814
rect 430 49698 59570 49814
rect 9 49142 59631 49698
rect 9 49026 70 49142
rect 430 49026 59570 49142
rect 9 48470 59631 49026
rect 9 48354 70 48470
rect 430 48354 59570 48470
rect 9 47798 59631 48354
rect 9 47682 70 47798
rect 430 47682 59570 47798
rect 9 47462 59631 47682
rect 9 47346 70 47462
rect 430 47346 59570 47462
rect 9 46790 59631 47346
rect 9 46674 70 46790
rect 430 46674 59570 46790
rect 9 46118 59631 46674
rect 9 46002 70 46118
rect 430 46002 59570 46118
rect 9 45446 59631 46002
rect 9 45330 70 45446
rect 430 45330 59570 45446
rect 9 45110 59631 45330
rect 9 44994 70 45110
rect 430 44994 59570 45110
rect 9 44438 59631 44994
rect 9 44322 70 44438
rect 430 44322 59570 44438
rect 9 43766 59631 44322
rect 9 43650 70 43766
rect 430 43650 59570 43766
rect 9 43430 59631 43650
rect 9 43314 70 43430
rect 430 43314 59570 43430
rect 9 42758 59631 43314
rect 9 42642 70 42758
rect 430 42642 59570 42758
rect 9 42086 59631 42642
rect 9 41970 70 42086
rect 430 41970 59570 42086
rect 9 41414 59631 41970
rect 9 41298 70 41414
rect 430 41298 59570 41414
rect 9 41078 59631 41298
rect 9 40962 70 41078
rect 430 40962 59570 41078
rect 9 40406 59631 40962
rect 9 40290 70 40406
rect 430 40290 59570 40406
rect 9 39734 59631 40290
rect 9 39618 70 39734
rect 430 39618 59570 39734
rect 9 39398 59631 39618
rect 9 39282 70 39398
rect 430 39282 59570 39398
rect 9 38726 59631 39282
rect 9 38610 70 38726
rect 430 38610 59570 38726
rect 9 38054 59631 38610
rect 9 37938 70 38054
rect 430 37938 59570 38054
rect 9 37382 59631 37938
rect 9 37266 70 37382
rect 430 37266 59570 37382
rect 9 37046 59631 37266
rect 9 36930 70 37046
rect 430 36930 59570 37046
rect 9 36374 59631 36930
rect 9 36258 70 36374
rect 430 36258 59570 36374
rect 9 35702 59631 36258
rect 9 35586 70 35702
rect 430 35586 59570 35702
rect 9 35030 59631 35586
rect 9 34914 70 35030
rect 430 34914 59570 35030
rect 9 34694 59631 34914
rect 9 34578 70 34694
rect 430 34578 59570 34694
rect 9 34022 59631 34578
rect 9 33906 70 34022
rect 430 33906 59570 34022
rect 9 33350 59631 33906
rect 9 33234 70 33350
rect 430 33234 59570 33350
rect 9 33014 59631 33234
rect 9 32898 70 33014
rect 430 32898 59570 33014
rect 9 32342 59631 32898
rect 9 32226 70 32342
rect 430 32226 59570 32342
rect 9 31670 59631 32226
rect 9 31554 70 31670
rect 430 31554 59570 31670
rect 9 30998 59631 31554
rect 9 30882 70 30998
rect 430 30882 59570 30998
rect 9 30662 59631 30882
rect 9 30546 70 30662
rect 430 30546 59570 30662
rect 9 29990 59631 30546
rect 9 29874 70 29990
rect 430 29874 59570 29990
rect 9 29318 59631 29874
rect 9 29202 70 29318
rect 430 29202 59570 29318
rect 9 28982 59631 29202
rect 9 28866 70 28982
rect 430 28866 59570 28982
rect 9 28310 59631 28866
rect 9 28194 70 28310
rect 430 28194 59570 28310
rect 9 27638 59631 28194
rect 9 27522 70 27638
rect 430 27522 59570 27638
rect 9 26966 59631 27522
rect 9 26850 70 26966
rect 430 26850 59570 26966
rect 9 26630 59631 26850
rect 9 26514 70 26630
rect 430 26514 59570 26630
rect 9 25958 59631 26514
rect 9 25842 70 25958
rect 430 25842 59570 25958
rect 9 25286 59631 25842
rect 9 25170 70 25286
rect 430 25170 59570 25286
rect 9 24950 59631 25170
rect 9 24834 70 24950
rect 430 24834 59570 24950
rect 9 24278 59631 24834
rect 9 24162 70 24278
rect 430 24162 59570 24278
rect 9 23606 59631 24162
rect 9 23490 70 23606
rect 430 23490 59570 23606
rect 9 22934 59631 23490
rect 9 22818 70 22934
rect 430 22818 59570 22934
rect 9 22598 59631 22818
rect 9 22482 70 22598
rect 430 22482 59570 22598
rect 9 21926 59631 22482
rect 9 21810 70 21926
rect 430 21810 59570 21926
rect 9 21254 59631 21810
rect 9 21138 70 21254
rect 430 21138 59570 21254
rect 9 20582 59631 21138
rect 9 20466 70 20582
rect 430 20466 59570 20582
rect 9 20246 59631 20466
rect 9 20130 70 20246
rect 430 20130 59570 20246
rect 9 19574 59631 20130
rect 9 19458 70 19574
rect 430 19458 59570 19574
rect 9 18902 59631 19458
rect 9 18786 70 18902
rect 430 18786 59570 18902
rect 9 18566 59631 18786
rect 9 18450 70 18566
rect 430 18450 59570 18566
rect 9 17894 59631 18450
rect 9 17778 70 17894
rect 430 17778 59570 17894
rect 9 17222 59631 17778
rect 9 17106 70 17222
rect 430 17106 59570 17222
rect 9 16550 59631 17106
rect 9 16434 70 16550
rect 430 16434 59570 16550
rect 9 16214 59631 16434
rect 9 16098 70 16214
rect 430 16098 59570 16214
rect 9 15542 59631 16098
rect 9 15426 70 15542
rect 430 15426 59570 15542
rect 9 14870 59631 15426
rect 9 14754 70 14870
rect 430 14754 59570 14870
rect 9 14534 59631 14754
rect 9 14418 70 14534
rect 430 14418 59570 14534
rect 9 13862 59631 14418
rect 9 13746 70 13862
rect 430 13746 59570 13862
rect 9 13190 59631 13746
rect 9 13074 70 13190
rect 430 13074 59570 13190
rect 9 12518 59631 13074
rect 9 12402 70 12518
rect 430 12402 59570 12518
rect 9 12182 59631 12402
rect 9 12066 70 12182
rect 430 12066 59570 12182
rect 9 11510 59631 12066
rect 9 11394 70 11510
rect 430 11394 59570 11510
rect 9 10838 59631 11394
rect 9 10722 70 10838
rect 430 10722 59570 10838
rect 9 10166 59631 10722
rect 9 10050 70 10166
rect 430 10050 59570 10166
rect 9 9830 59631 10050
rect 9 9714 70 9830
rect 430 9714 59570 9830
rect 9 9158 59631 9714
rect 9 9042 70 9158
rect 430 9042 59570 9158
rect 9 8486 59631 9042
rect 9 8370 70 8486
rect 430 8370 59570 8486
rect 9 8150 59631 8370
rect 9 8034 70 8150
rect 430 8034 59570 8150
rect 9 7478 59631 8034
rect 9 7362 70 7478
rect 430 7362 59570 7478
rect 9 6806 59631 7362
rect 9 6690 70 6806
rect 430 6690 59570 6806
rect 9 6134 59631 6690
rect 9 6018 70 6134
rect 430 6018 59570 6134
rect 9 5798 59631 6018
rect 9 5682 70 5798
rect 430 5682 59570 5798
rect 9 5126 59631 5682
rect 9 5010 70 5126
rect 430 5010 59570 5126
rect 9 4454 59631 5010
rect 9 4338 70 4454
rect 430 4338 59570 4454
rect 9 4118 59631 4338
rect 9 4002 70 4118
rect 430 4002 59570 4118
rect 9 3446 59631 4002
rect 9 3330 70 3446
rect 430 3330 59570 3446
rect 9 2774 59631 3330
rect 9 2658 70 2774
rect 430 2658 59570 2774
rect 9 2102 59631 2658
rect 9 1986 70 2102
rect 430 1986 59570 2102
rect 9 1766 59631 1986
rect 9 1650 70 1766
rect 430 1650 59570 1766
rect 9 1094 59631 1650
rect 9 978 70 1094
rect 430 978 59570 1094
rect 9 798 59631 978
<< metal4 >>
rect 2224 1538 2384 58438
rect 9904 1538 10064 58438
rect 17584 1538 17744 58438
rect 25264 1538 25424 58438
rect 32944 1538 33104 58438
rect 40624 1538 40784 58438
rect 48304 1538 48464 58438
rect 55984 1538 56144 58438
<< obsm4 >>
rect 1582 1508 2194 53975
rect 2414 1508 9874 53975
rect 10094 1508 17554 53975
rect 17774 1508 25234 53975
rect 25454 1508 32914 53975
rect 33134 1508 40594 53975
rect 40814 1508 48274 53975
rect 48494 1508 55954 53975
rect 56174 1508 59178 53975
rect 1582 1465 59178 1508
<< labels >>
rlabel metal3 s 100 41328 400 41384 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 100 42000 400 42056 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 100 20496 400 20552 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 100 36288 400 36344 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 100 24864 400 24920 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 100 21168 400 21224 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 31584 59600 31640 59900 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 59600 12096 59900 12152 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 59600 56448 59900 56504 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 40320 59600 40376 59900 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 58800 100 58856 400 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 7392 59600 7448 59900 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 47712 59600 47768 59900 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 42000 100 42056 400 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 59808 59600 59864 59900 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 59600 51744 59900 51800 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 49728 100 49784 400 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 8064 100 8120 400 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 100 50064 400 50120 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 100 40992 400 41048 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 100 46704 400 46760 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 100 37296 400 37352 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 59600 59472 59900 59528 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 39312 100 39368 400 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 100 25200 400 25256 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 50736 100 50792 400 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 100 6048 400 6104 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 100 53760 400 53816 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 53760 59600 53816 59900 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 59600 53088 59900 53144 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 59600 45360 59900 45416 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 59600 58800 59900 58856 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 59600 26880 59900 26936 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 100 11424 400 11480 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 59600 11424 59900 11480 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 49056 59600 49112 59900 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 100 27552 400 27608 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 100 30912 400 30968 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 59600 42000 59900 42056 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 59600 38640 59900 38696 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 2016 59600 2072 59900 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 36960 100 37016 400 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 100 15456 400 15512 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 54768 100 54824 400 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 37968 59600 38024 59900 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 17136 100 17192 400 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 5712 100 5768 400 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 2688 59600 2744 59900 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 21168 59600 21224 59900 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 16128 59600 16184 59900 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 34608 59600 34664 59900 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 51408 100 51464 400 6 io_oeb[21]
port 52 nsew signal output
rlabel metal3 s 59600 15456 59900 15512 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 58128 59600 58184 59900 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 100 17136 400 17192 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 100 8400 400 8456 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 100 54768 400 54824 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 50064 100 50120 400 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 1008 59600 1064 59900 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 59600 30576 59900 30632 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 59600 22848 59900 22904 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 56448 100 56504 400 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 100 18480 400 18536 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 52416 59600 52472 59900 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 59600 9744 59900 9800 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 100 49056 400 49112 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 59600 54096 59900 54152 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 33264 59600 33320 59900 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 59600 24192 59900 24248 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 100 45024 400 45080 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 100 8064 400 8120 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 43680 59600 43736 59900 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 100 47376 400 47432 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 28896 59600 28952 59900 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 100 29904 400 29960 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 59600 58128 59900 58184 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 9744 59600 9800 59900 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 18480 59600 18536 59900 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 38640 100 38696 400 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 58800 59600 58856 59900 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 100 59808 400 59864 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 100 44352 400 44408 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 24192 100 24248 400 6 io_out[15]
port 83 nsew signal output
rlabel metal3 s 59600 50064 59900 50120 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 6720 100 6776 400 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 55776 100 55832 400 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 13104 59600 13160 59900 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 4032 100 4088 400 6 io_out[1]
port 88 nsew signal output
rlabel metal3 s 59600 5712 59900 5768 6 io_out[20]
port 89 nsew signal output
rlabel metal3 s 100 39648 400 39704 6 io_out[21]
port 90 nsew signal output
rlabel metal3 s 59600 13104 59900 13160 6 io_out[22]
port 91 nsew signal output
rlabel metal3 s 100 22512 400 22568 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 52416 100 52472 400 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 59600 1680 59900 1736 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 25200 100 25256 400 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 20160 100 20216 400 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 42000 59600 42056 59900 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 40992 100 41048 400 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 59600 21168 59900 21224 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 54768 59600 54824 59900 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 21168 100 21224 400 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 37296 59600 37352 59900 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 100 21840 400 21896 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 39648 100 39704 400 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 35616 100 35672 400 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 14448 100 14504 400 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 100 2688 400 2744 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 27552 59600 27608 59900 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 27552 100 27608 400 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 25200 59600 25256 59900 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 100 10752 400 10808 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 100 33936 400 33992 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 43680 100 43736 400 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 15456 100 15512 400 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 100 30576 400 30632 6 la_data_in[0]
port 115 nsew signal input
rlabel metal3 s 59600 55776 59900 55832 6 la_data_in[10]
port 116 nsew signal input
rlabel metal3 s 59600 26544 59900 26600 6 la_data_in[11]
port 117 nsew signal input
rlabel metal2 s 18480 100 18536 400 6 la_data_in[12]
port 118 nsew signal input
rlabel metal2 s 24192 59600 24248 59900 6 la_data_in[13]
port 119 nsew signal input
rlabel metal3 s 100 52416 400 52472 6 la_data_in[14]
port 120 nsew signal input
rlabel metal3 s 59600 43344 59900 43400 6 la_data_in[15]
port 121 nsew signal input
rlabel metal2 s 5712 59600 5768 59900 6 la_data_in[16]
port 122 nsew signal input
rlabel metal3 s 59600 9072 59900 9128 6 la_data_in[17]
port 123 nsew signal input
rlabel metal2 s 29904 59600 29960 59900 6 la_data_in[18]
port 124 nsew signal input
rlabel metal3 s 100 9072 400 9128 6 la_data_in[19]
port 125 nsew signal input
rlabel metal2 s 13776 59600 13832 59900 6 la_data_in[1]
port 126 nsew signal input
rlabel metal3 s 59600 12432 59900 12488 6 la_data_in[20]
port 127 nsew signal input
rlabel metal3 s 100 45360 400 45416 6 la_data_in[21]
port 128 nsew signal input
rlabel metal3 s 100 26544 400 26600 6 la_data_in[22]
port 129 nsew signal input
rlabel metal3 s 59600 45024 59900 45080 6 la_data_in[23]
port 130 nsew signal input
rlabel metal2 s 30576 59600 30632 59900 6 la_data_in[24]
port 131 nsew signal input
rlabel metal2 s 12432 59600 12488 59900 6 la_data_in[25]
port 132 nsew signal input
rlabel metal2 s 36960 59600 37016 59900 6 la_data_in[26]
port 133 nsew signal input
rlabel metal3 s 100 54096 400 54152 6 la_data_in[27]
port 134 nsew signal input
rlabel metal3 s 100 56448 400 56504 6 la_data_in[28]
port 135 nsew signal input
rlabel metal3 s 59600 14784 59900 14840 6 la_data_in[29]
port 136 nsew signal input
rlabel metal2 s 26544 59600 26600 59900 6 la_data_in[2]
port 137 nsew signal input
rlabel metal3 s 100 4368 400 4424 6 la_data_in[30]
port 138 nsew signal input
rlabel metal2 s 50736 59600 50792 59900 6 la_data_in[31]
port 139 nsew signal input
rlabel metal3 s 100 24192 400 24248 6 la_data_in[32]
port 140 nsew signal input
rlabel metal3 s 100 40320 400 40376 6 la_data_in[33]
port 141 nsew signal input
rlabel metal2 s 4368 59600 4424 59900 6 la_data_in[34]
port 142 nsew signal input
rlabel metal3 s 100 53088 400 53144 6 la_data_in[35]
port 143 nsew signal input
rlabel metal2 s 42672 100 42728 400 6 la_data_in[36]
port 144 nsew signal input
rlabel metal3 s 100 58800 400 58856 6 la_data_in[37]
port 145 nsew signal input
rlabel metal2 s 26880 100 26936 400 6 la_data_in[38]
port 146 nsew signal input
rlabel metal2 s 32928 59600 32984 59900 6 la_data_in[39]
port 147 nsew signal input
rlabel metal3 s 59600 32928 59900 32984 6 la_data_in[3]
port 148 nsew signal input
rlabel metal2 s 20496 100 20552 400 6 la_data_in[40]
port 149 nsew signal input
rlabel metal2 s 28896 100 28952 400 6 la_data_in[41]
port 150 nsew signal input
rlabel metal3 s 100 20160 400 20216 6 la_data_in[42]
port 151 nsew signal input
rlabel metal2 s 56448 59600 56504 59900 6 la_data_in[43]
port 152 nsew signal input
rlabel metal3 s 59600 336 59900 392 6 la_data_in[44]
port 153 nsew signal input
rlabel metal2 s 19488 100 19544 400 6 la_data_in[45]
port 154 nsew signal input
rlabel metal3 s 59600 43680 59900 43736 6 la_data_in[46]
port 155 nsew signal input
rlabel metal2 s 37296 100 37352 400 6 la_data_in[47]
port 156 nsew signal input
rlabel metal2 s 28224 59600 28280 59900 6 la_data_in[48]
port 157 nsew signal input
rlabel metal2 s 22848 59600 22904 59900 6 la_data_in[49]
port 158 nsew signal input
rlabel metal2 s 5040 59600 5096 59900 6 la_data_in[4]
port 159 nsew signal input
rlabel metal2 s 23520 59600 23576 59900 6 la_data_in[50]
port 160 nsew signal input
rlabel metal2 s 28224 100 28280 400 6 la_data_in[51]
port 161 nsew signal input
rlabel metal3 s 59600 20160 59900 20216 6 la_data_in[52]
port 162 nsew signal input
rlabel metal2 s 46704 59600 46760 59900 6 la_data_in[53]
port 163 nsew signal input
rlabel metal2 s 42672 59600 42728 59900 6 la_data_in[54]
port 164 nsew signal input
rlabel metal3 s 100 16128 400 16184 6 la_data_in[55]
port 165 nsew signal input
rlabel metal3 s 100 17808 400 17864 6 la_data_in[56]
port 166 nsew signal input
rlabel metal2 s 1680 59600 1736 59900 6 la_data_in[57]
port 167 nsew signal input
rlabel metal2 s 21840 100 21896 400 6 la_data_in[58]
port 168 nsew signal input
rlabel metal3 s 59600 54768 59900 54824 6 la_data_in[59]
port 169 nsew signal input
rlabel metal2 s 10080 100 10136 400 6 la_data_in[5]
port 170 nsew signal input
rlabel metal3 s 59600 39648 59900 39704 6 la_data_in[60]
port 171 nsew signal input
rlabel metal3 s 100 1680 400 1736 6 la_data_in[61]
port 172 nsew signal input
rlabel metal2 s 34944 100 35000 400 6 la_data_in[62]
port 173 nsew signal input
rlabel metal2 s 15456 59600 15512 59900 6 la_data_in[63]
port 174 nsew signal input
rlabel metal2 s 12096 100 12152 400 6 la_data_in[6]
port 175 nsew signal input
rlabel metal3 s 59600 21840 59900 21896 6 la_data_in[7]
port 176 nsew signal input
rlabel metal3 s 100 1008 400 1064 6 la_data_in[8]
port 177 nsew signal input
rlabel metal2 s 54096 59600 54152 59900 6 la_data_in[9]
port 178 nsew signal input
rlabel metal2 s 51744 59600 51800 59900 6 la_data_out[0]
port 179 nsew signal output
rlabel metal3 s 59600 32256 59900 32312 6 la_data_out[10]
port 180 nsew signal output
rlabel metal3 s 100 2016 400 2072 6 la_data_out[11]
port 181 nsew signal output
rlabel metal3 s 100 43344 400 43400 6 la_data_out[12]
port 182 nsew signal output
rlabel metal2 s 22512 100 22568 400 6 la_data_out[13]
port 183 nsew signal output
rlabel metal3 s 59600 24864 59900 24920 6 la_data_out[14]
port 184 nsew signal output
rlabel metal3 s 100 51408 400 51464 6 la_data_out[15]
port 185 nsew signal output
rlabel metal3 s 59600 33264 59900 33320 6 la_data_out[16]
port 186 nsew signal output
rlabel metal2 s 29232 59600 29288 59900 6 la_data_out[17]
port 187 nsew signal output
rlabel metal3 s 59600 49728 59900 49784 6 la_data_out[18]
port 188 nsew signal output
rlabel metal2 s 31584 100 31640 400 6 la_data_out[19]
port 189 nsew signal output
rlabel metal3 s 59600 28224 59900 28280 6 la_data_out[1]
port 190 nsew signal output
rlabel metal3 s 59600 8400 59900 8456 6 la_data_out[20]
port 191 nsew signal output
rlabel metal3 s 100 59472 400 59528 6 la_data_out[21]
port 192 nsew signal output
rlabel metal3 s 59600 37296 59900 37352 6 la_data_out[22]
port 193 nsew signal output
rlabel metal2 s 17808 100 17864 400 6 la_data_out[23]
port 194 nsew signal output
rlabel metal3 s 100 26880 400 26936 6 la_data_out[24]
port 195 nsew signal output
rlabel metal2 s 32256 100 32312 400 6 la_data_out[25]
port 196 nsew signal output
rlabel metal3 s 100 58128 400 58184 6 la_data_out[26]
port 197 nsew signal output
rlabel metal2 s 36288 59600 36344 59900 6 la_data_out[27]
port 198 nsew signal output
rlabel metal3 s 59600 47712 59900 47768 6 la_data_out[28]
port 199 nsew signal output
rlabel metal2 s 25872 100 25928 400 6 la_data_out[29]
port 200 nsew signal output
rlabel metal3 s 100 13776 400 13832 6 la_data_out[2]
port 201 nsew signal output
rlabel metal3 s 59600 27552 59900 27608 6 la_data_out[30]
port 202 nsew signal output
rlabel metal3 s 59600 2688 59900 2744 6 la_data_out[31]
port 203 nsew signal output
rlabel metal2 s 34944 59600 35000 59900 6 la_data_out[32]
port 204 nsew signal output
rlabel metal3 s 59600 10752 59900 10808 6 la_data_out[33]
port 205 nsew signal output
rlabel metal2 s 29232 100 29288 400 6 la_data_out[34]
port 206 nsew signal output
rlabel metal2 s 32256 59600 32312 59900 6 la_data_out[35]
port 207 nsew signal output
rlabel metal3 s 59600 48384 59900 48440 6 la_data_out[36]
port 208 nsew signal output
rlabel metal3 s 59600 23520 59900 23576 6 la_data_out[37]
port 209 nsew signal output
rlabel metal3 s 59600 1008 59900 1064 6 la_data_out[38]
port 210 nsew signal output
rlabel metal3 s 59600 8064 59900 8120 6 la_data_out[39]
port 211 nsew signal output
rlabel metal3 s 100 9744 400 9800 6 la_data_out[3]
port 212 nsew signal output
rlabel metal2 s 58128 100 58184 400 6 la_data_out[40]
port 213 nsew signal output
rlabel metal3 s 59600 18480 59900 18536 6 la_data_out[41]
port 214 nsew signal output
rlabel metal3 s 59600 50736 59900 50792 6 la_data_out[42]
port 215 nsew signal output
rlabel metal2 s 3360 100 3416 400 6 la_data_out[43]
port 216 nsew signal output
rlabel metal2 s 24864 100 24920 400 6 la_data_out[44]
port 217 nsew signal output
rlabel metal2 s 9072 59600 9128 59900 6 la_data_out[45]
port 218 nsew signal output
rlabel metal2 s 8400 59600 8456 59900 6 la_data_out[46]
port 219 nsew signal output
rlabel metal3 s 100 42672 400 42728 6 la_data_out[47]
port 220 nsew signal output
rlabel metal2 s 13776 100 13832 400 6 la_data_out[48]
port 221 nsew signal output
rlabel metal2 s 54096 100 54152 400 6 la_data_out[49]
port 222 nsew signal output
rlabel metal2 s 33936 59600 33992 59900 6 la_data_out[4]
port 223 nsew signal output
rlabel metal2 s 20496 59600 20552 59900 6 la_data_out[50]
port 224 nsew signal output
rlabel metal3 s 100 57792 400 57848 6 la_data_out[51]
port 225 nsew signal output
rlabel metal3 s 59600 4032 59900 4088 6 la_data_out[52]
port 226 nsew signal output
rlabel metal3 s 100 57120 400 57176 6 la_data_out[53]
port 227 nsew signal output
rlabel metal3 s 59600 40992 59900 41048 6 la_data_out[54]
port 228 nsew signal output
rlabel metal2 s 22512 59600 22568 59900 6 la_data_out[55]
port 229 nsew signal output
rlabel metal3 s 59600 14448 59900 14504 6 la_data_out[56]
port 230 nsew signal output
rlabel metal2 s 45360 59600 45416 59900 6 la_data_out[57]
port 231 nsew signal output
rlabel metal3 s 59600 41328 59900 41384 6 la_data_out[58]
port 232 nsew signal output
rlabel metal3 s 100 22848 400 22904 6 la_data_out[59]
port 233 nsew signal output
rlabel metal3 s 59600 35616 59900 35672 6 la_data_out[5]
port 234 nsew signal output
rlabel metal2 s 48384 59600 48440 59900 6 la_data_out[60]
port 235 nsew signal output
rlabel metal2 s 16128 100 16184 400 6 la_data_out[61]
port 236 nsew signal output
rlabel metal2 s 51744 100 51800 400 6 la_data_out[62]
port 237 nsew signal output
rlabel metal3 s 59600 4368 59900 4424 6 la_data_out[63]
port 238 nsew signal output
rlabel metal3 s 59600 17136 59900 17192 6 la_data_out[6]
port 239 nsew signal output
rlabel metal2 s 57792 59600 57848 59900 6 la_data_out[7]
port 240 nsew signal output
rlabel metal3 s 100 3360 400 3416 6 la_data_out[8]
port 241 nsew signal output
rlabel metal3 s 59600 28896 59900 28952 6 la_data_out[9]
port 242 nsew signal output
rlabel metal3 s 59600 22512 59900 22568 6 la_oenb[0]
port 243 nsew signal input
rlabel metal3 s 59600 42672 59900 42728 6 la_oenb[10]
port 244 nsew signal input
rlabel metal3 s 59600 33936 59900 33992 6 la_oenb[11]
port 245 nsew signal input
rlabel metal2 s 336 59600 392 59900 6 la_oenb[12]
port 246 nsew signal input
rlabel metal3 s 100 47712 400 47768 6 la_oenb[13]
port 247 nsew signal input
rlabel metal2 s 44352 100 44408 400 6 la_oenb[14]
port 248 nsew signal input
rlabel metal2 s 53088 100 53144 400 6 la_oenb[15]
port 249 nsew signal input
rlabel metal2 s 8400 100 8456 400 6 la_oenb[16]
port 250 nsew signal input
rlabel metal3 s 100 7392 400 7448 6 la_oenb[17]
port 251 nsew signal input
rlabel metal2 s 4032 59600 4088 59900 6 la_oenb[18]
port 252 nsew signal input
rlabel metal3 s 59600 5040 59900 5096 6 la_oenb[19]
port 253 nsew signal input
rlabel metal2 s 11424 59600 11480 59900 6 la_oenb[1]
port 254 nsew signal input
rlabel metal3 s 100 34944 400 35000 6 la_oenb[20]
port 255 nsew signal input
rlabel metal2 s 24864 59600 24920 59900 6 la_oenb[21]
port 256 nsew signal input
rlabel metal2 s 44352 59600 44408 59900 6 la_oenb[22]
port 257 nsew signal input
rlabel metal2 s 16464 100 16520 400 6 la_oenb[23]
port 258 nsew signal input
rlabel metal3 s 59600 36960 59900 37016 6 la_oenb[24]
port 259 nsew signal input
rlabel metal2 s 53760 100 53816 400 6 la_oenb[25]
port 260 nsew signal input
rlabel metal2 s 12096 59600 12152 59900 6 la_oenb[26]
port 261 nsew signal input
rlabel metal2 s 10752 100 10808 400 6 la_oenb[27]
port 262 nsew signal input
rlabel metal3 s 100 36960 400 37016 6 la_oenb[28]
port 263 nsew signal input
rlabel metal3 s 59600 57120 59900 57176 6 la_oenb[29]
port 264 nsew signal input
rlabel metal2 s 59472 59600 59528 59900 6 la_oenb[2]
port 265 nsew signal input
rlabel metal3 s 59600 51408 59900 51464 6 la_oenb[30]
port 266 nsew signal input
rlabel metal2 s 25872 59600 25928 59900 6 la_oenb[31]
port 267 nsew signal input
rlabel metal3 s 59600 49056 59900 49112 6 la_oenb[32]
port 268 nsew signal input
rlabel metal2 s 30576 100 30632 400 6 la_oenb[33]
port 269 nsew signal input
rlabel metal2 s 10080 59600 10136 59900 6 la_oenb[34]
port 270 nsew signal input
rlabel metal2 s 1680 100 1736 400 6 la_oenb[35]
port 271 nsew signal input
rlabel metal2 s 336 100 392 400 6 la_oenb[36]
port 272 nsew signal input
rlabel metal2 s 8064 59600 8120 59900 6 la_oenb[37]
port 273 nsew signal input
rlabel metal2 s 30912 100 30968 400 6 la_oenb[38]
port 274 nsew signal input
rlabel metal3 s 100 25872 400 25928 6 la_oenb[39]
port 275 nsew signal input
rlabel metal3 s 100 32928 400 32984 6 la_oenb[3]
port 276 nsew signal input
rlabel metal3 s 59600 7392 59900 7448 6 la_oenb[40]
port 277 nsew signal input
rlabel metal2 s 21840 59600 21896 59900 6 la_oenb[41]
port 278 nsew signal input
rlabel metal3 s 100 37968 400 38024 6 la_oenb[42]
port 279 nsew signal input
rlabel metal2 s 11424 100 11480 400 6 la_oenb[43]
port 280 nsew signal input
rlabel metal2 s 26544 100 26600 400 6 la_oenb[44]
port 281 nsew signal input
rlabel metal2 s 49728 59600 49784 59900 6 la_oenb[45]
port 282 nsew signal input
rlabel metal2 s 47712 100 47768 400 6 la_oenb[46]
port 283 nsew signal input
rlabel metal3 s 100 6720 400 6776 6 la_oenb[47]
port 284 nsew signal input
rlabel metal3 s 100 43680 400 43736 6 la_oenb[48]
port 285 nsew signal input
rlabel metal3 s 100 336 400 392 6 la_oenb[49]
port 286 nsew signal input
rlabel metal3 s 100 55776 400 55832 6 la_oenb[4]
port 287 nsew signal input
rlabel metal2 s 46032 100 46088 400 6 la_oenb[50]
port 288 nsew signal input
rlabel metal2 s 19488 59600 19544 59900 6 la_oenb[51]
port 289 nsew signal input
rlabel metal2 s 59472 100 59528 400 6 la_oenb[52]
port 290 nsew signal input
rlabel metal3 s 59600 37968 59900 38024 6 la_oenb[53]
port 291 nsew signal input
rlabel metal3 s 100 32256 400 32312 6 la_oenb[54]
port 292 nsew signal input
rlabel metal3 s 59600 30912 59900 30968 6 la_oenb[55]
port 293 nsew signal input
rlabel metal2 s 45360 100 45416 400 6 la_oenb[56]
port 294 nsew signal input
rlabel metal2 s 53088 59600 53144 59900 6 la_oenb[57]
port 295 nsew signal input
rlabel metal3 s 59600 6048 59900 6104 6 la_oenb[58]
port 296 nsew signal input
rlabel metal2 s 35616 59600 35672 59900 6 la_oenb[59]
port 297 nsew signal input
rlabel metal2 s 55440 100 55496 400 6 la_oenb[5]
port 298 nsew signal input
rlabel metal3 s 100 29232 400 29288 6 la_oenb[60]
port 299 nsew signal input
rlabel metal2 s 7392 100 7448 400 6 la_oenb[61]
port 300 nsew signal input
rlabel metal3 s 59600 29904 59900 29960 6 la_oenb[62]
port 301 nsew signal input
rlabel metal3 s 100 14448 400 14504 6 la_oenb[63]
port 302 nsew signal input
rlabel metal3 s 59600 39312 59900 39368 6 la_oenb[6]
port 303 nsew signal input
rlabel metal2 s 14784 100 14840 400 6 la_oenb[7]
port 304 nsew signal input
rlabel metal2 s 57120 100 57176 400 6 la_oenb[8]
port 305 nsew signal input
rlabel metal2 s 17136 59600 17192 59900 6 la_oenb[9]
port 306 nsew signal input
rlabel metal2 s 51408 59600 51464 59900 6 user_clock2
port 307 nsew signal input
rlabel metal3 s 59600 46032 59900 46088 6 user_irq[0]
port 308 nsew signal output
rlabel metal2 s 14784 59600 14840 59900 6 user_irq[1]
port 309 nsew signal output
rlabel metal3 s 100 38640 400 38696 6 user_irq[2]
port 310 nsew signal output
rlabel metal4 s 2224 1538 2384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal3 s 59600 10080 59900 10136 6 wb_clk_i
port 313 nsew signal input
rlabel metal2 s 10752 59600 10808 59900 6 wb_rst_i
port 314 nsew signal input
rlabel metal3 s 59600 20496 59900 20552 6 wbs_ack_o
port 315 nsew signal output
rlabel metal2 s 39648 59600 39704 59900 6 wbs_adr_i[0]
port 316 nsew signal input
rlabel metal2 s 26880 59600 26936 59900 6 wbs_adr_i[10]
port 317 nsew signal input
rlabel metal3 s 100 34608 400 34664 6 wbs_adr_i[11]
port 318 nsew signal input
rlabel metal2 s 5040 100 5096 400 6 wbs_adr_i[12]
port 319 nsew signal input
rlabel metal2 s 33264 100 33320 400 6 wbs_adr_i[13]
port 320 nsew signal input
rlabel metal3 s 100 5712 400 5768 6 wbs_adr_i[14]
port 321 nsew signal input
rlabel metal3 s 59600 40320 59900 40376 6 wbs_adr_i[15]
port 322 nsew signal input
rlabel metal2 s 37968 100 38024 400 6 wbs_adr_i[16]
port 323 nsew signal input
rlabel metal3 s 100 33264 400 33320 6 wbs_adr_i[17]
port 324 nsew signal input
rlabel metal3 s 59600 18816 59900 18872 6 wbs_adr_i[18]
port 325 nsew signal input
rlabel metal2 s 57792 100 57848 400 6 wbs_adr_i[19]
port 326 nsew signal input
rlabel metal3 s 100 4032 400 4088 6 wbs_adr_i[1]
port 327 nsew signal input
rlabel metal2 s 55776 59600 55832 59900 6 wbs_adr_i[20]
port 328 nsew signal input
rlabel metal2 s 33936 100 33992 400 6 wbs_adr_i[21]
port 329 nsew signal input
rlabel metal2 s 48384 100 48440 400 6 wbs_adr_i[22]
port 330 nsew signal input
rlabel metal3 s 59600 13776 59900 13832 6 wbs_adr_i[23]
port 331 nsew signal input
rlabel metal2 s 6720 59600 6776 59900 6 wbs_adr_i[24]
port 332 nsew signal input
rlabel metal3 s 100 10080 400 10136 6 wbs_adr_i[25]
port 333 nsew signal input
rlabel metal2 s 6048 100 6104 400 6 wbs_adr_i[26]
port 334 nsew signal input
rlabel metal2 s 20160 59600 20216 59900 6 wbs_adr_i[27]
port 335 nsew signal input
rlabel metal3 s 59600 34944 59900 35000 6 wbs_adr_i[28]
port 336 nsew signal input
rlabel metal3 s 59600 57792 59900 57848 6 wbs_adr_i[29]
port 337 nsew signal input
rlabel metal2 s 23520 100 23576 400 6 wbs_adr_i[2]
port 338 nsew signal input
rlabel metal3 s 100 23520 400 23576 6 wbs_adr_i[30]
port 339 nsew signal input
rlabel metal3 s 59600 25200 59900 25256 6 wbs_adr_i[31]
port 340 nsew signal input
rlabel metal2 s 46704 100 46760 400 6 wbs_adr_i[3]
port 341 nsew signal input
rlabel metal2 s 46032 59600 46088 59900 6 wbs_adr_i[4]
port 342 nsew signal input
rlabel metal2 s 45024 100 45080 400 6 wbs_adr_i[5]
port 343 nsew signal input
rlabel metal3 s 100 14784 400 14840 6 wbs_adr_i[6]
port 344 nsew signal input
rlabel metal2 s 2688 100 2744 400 6 wbs_adr_i[7]
port 345 nsew signal input
rlabel metal3 s 59600 0 59900 56 6 wbs_adr_i[8]
port 346 nsew signal input
rlabel metal3 s 59600 16128 59900 16184 6 wbs_adr_i[9]
port 347 nsew signal input
rlabel metal2 s 18816 59600 18872 59900 6 wbs_cyc_i
port 348 nsew signal input
rlabel metal3 s 59600 52416 59900 52472 6 wbs_dat_i[0]
port 349 nsew signal input
rlabel metal3 s 100 46032 400 46088 6 wbs_dat_i[10]
port 350 nsew signal input
rlabel metal3 s 100 50736 400 50792 6 wbs_dat_i[11]
port 351 nsew signal input
rlabel metal3 s 100 48384 400 48440 6 wbs_dat_i[12]
port 352 nsew signal input
rlabel metal2 s 2016 100 2072 400 6 wbs_dat_i[13]
port 353 nsew signal input
rlabel metal3 s 100 12432 400 12488 6 wbs_dat_i[14]
port 354 nsew signal input
rlabel metal3 s 59600 31584 59900 31640 6 wbs_dat_i[15]
port 355 nsew signal input
rlabel metal2 s 34608 100 34664 400 6 wbs_dat_i[16]
port 356 nsew signal input
rlabel metal2 s 40992 59600 41048 59900 6 wbs_dat_i[17]
port 357 nsew signal input
rlabel metal2 s 55440 59600 55496 59900 6 wbs_dat_i[18]
port 358 nsew signal input
rlabel metal2 s 3360 59600 3416 59900 6 wbs_dat_i[19]
port 359 nsew signal input
rlabel metal2 s 9072 100 9128 400 6 wbs_dat_i[1]
port 360 nsew signal input
rlabel metal3 s 100 28224 400 28280 6 wbs_dat_i[20]
port 361 nsew signal input
rlabel metal2 s 57120 59600 57176 59900 6 wbs_dat_i[21]
port 362 nsew signal input
rlabel metal3 s 100 35616 400 35672 6 wbs_dat_i[22]
port 363 nsew signal input
rlabel metal3 s 59600 47376 59900 47432 6 wbs_dat_i[23]
port 364 nsew signal input
rlabel metal3 s 59600 19488 59900 19544 6 wbs_dat_i[24]
port 365 nsew signal input
rlabel metal2 s 41328 100 41384 400 6 wbs_dat_i[25]
port 366 nsew signal input
rlabel metal2 s 50064 59600 50120 59900 6 wbs_dat_i[26]
port 367 nsew signal input
rlabel metal2 s 14448 59600 14504 59900 6 wbs_dat_i[27]
port 368 nsew signal input
rlabel metal2 s 18816 100 18872 400 6 wbs_dat_i[28]
port 369 nsew signal input
rlabel metal3 s 59600 36288 59900 36344 6 wbs_dat_i[29]
port 370 nsew signal input
rlabel metal2 s 49056 100 49112 400 6 wbs_dat_i[2]
port 371 nsew signal input
rlabel metal3 s 59600 17808 59900 17864 6 wbs_dat_i[30]
port 372 nsew signal input
rlabel metal3 s 100 31584 400 31640 6 wbs_dat_i[31]
port 373 nsew signal input
rlabel metal3 s 59600 2016 59900 2072 6 wbs_dat_i[3]
port 374 nsew signal input
rlabel metal2 s 9744 100 9800 400 6 wbs_dat_i[4]
port 375 nsew signal input
rlabel metal2 s 29904 100 29960 400 6 wbs_dat_i[5]
port 376 nsew signal input
rlabel metal3 s 59600 25872 59900 25928 6 wbs_dat_i[6]
port 377 nsew signal input
rlabel metal2 s 47376 59600 47432 59900 6 wbs_dat_i[7]
port 378 nsew signal input
rlabel metal3 s 59600 53760 59900 53816 6 wbs_dat_i[8]
port 379 nsew signal input
rlabel metal3 s 59600 3360 59900 3416 6 wbs_dat_i[9]
port 380 nsew signal input
rlabel metal3 s 100 12096 400 12152 6 wbs_dat_o[0]
port 381 nsew signal output
rlabel metal3 s 59600 34608 59900 34664 6 wbs_dat_o[10]
port 382 nsew signal output
rlabel metal2 s 1008 100 1064 400 6 wbs_dat_o[11]
port 383 nsew signal output
rlabel metal3 s 59600 55440 59900 55496 6 wbs_dat_o[12]
port 384 nsew signal output
rlabel metal2 s 45024 59600 45080 59900 6 wbs_dat_o[13]
port 385 nsew signal output
rlabel metal3 s 59600 6720 59900 6776 6 wbs_dat_o[14]
port 386 nsew signal output
rlabel metal2 s 43344 59600 43400 59900 6 wbs_dat_o[15]
port 387 nsew signal output
rlabel metal3 s 100 16464 400 16520 6 wbs_dat_o[16]
port 388 nsew signal output
rlabel metal3 s 100 18816 400 18872 6 wbs_dat_o[17]
port 389 nsew signal output
rlabel metal2 s 40320 100 40376 400 6 wbs_dat_o[18]
port 390 nsew signal output
rlabel metal2 s 0 100 56 400 6 wbs_dat_o[19]
port 391 nsew signal output
rlabel metal2 s 47376 100 47432 400 6 wbs_dat_o[1]
port 392 nsew signal output
rlabel metal3 s 100 28896 400 28952 6 wbs_dat_o[20]
port 393 nsew signal output
rlabel metal3 s 100 51744 400 51800 6 wbs_dat_o[21]
port 394 nsew signal output
rlabel metal2 s 16464 59600 16520 59900 6 wbs_dat_o[22]
port 395 nsew signal output
rlabel metal3 s 100 19488 400 19544 6 wbs_dat_o[23]
port 396 nsew signal output
rlabel metal2 s 12432 100 12488 400 6 wbs_dat_o[24]
port 397 nsew signal output
rlabel metal2 s 4368 100 4424 400 6 wbs_dat_o[25]
port 398 nsew signal output
rlabel metal2 s 30912 59600 30968 59900 6 wbs_dat_o[26]
port 399 nsew signal output
rlabel metal2 s 17808 59600 17864 59900 6 wbs_dat_o[27]
port 400 nsew signal output
rlabel metal2 s 32928 100 32984 400 6 wbs_dat_o[28]
port 401 nsew signal output
rlabel metal2 s 41328 59600 41384 59900 6 wbs_dat_o[29]
port 402 nsew signal output
rlabel metal3 s 59600 16464 59900 16520 6 wbs_dat_o[2]
port 403 nsew signal output
rlabel metal3 s 100 39312 400 39368 6 wbs_dat_o[30]
port 404 nsew signal output
rlabel metal3 s 59600 46704 59900 46760 6 wbs_dat_o[31]
port 405 nsew signal output
rlabel metal2 s 13104 100 13160 400 6 wbs_dat_o[3]
port 406 nsew signal output
rlabel metal2 s 22848 100 22904 400 6 wbs_dat_o[4]
port 407 nsew signal output
rlabel metal3 s 100 5040 400 5096 6 wbs_dat_o[5]
port 408 nsew signal output
rlabel metal3 s 59600 44352 59900 44408 6 wbs_dat_o[6]
port 409 nsew signal output
rlabel metal2 s 36288 100 36344 400 6 wbs_dat_o[7]
port 410 nsew signal output
rlabel metal2 s 39312 59600 39368 59900 6 wbs_dat_o[8]
port 411 nsew signal output
rlabel metal2 s 38640 59600 38696 59900 6 wbs_dat_o[9]
port 412 nsew signal output
rlabel metal3 s 100 55440 400 55496 6 wbs_sel_i[0]
port 413 nsew signal input
rlabel metal2 s 6048 59600 6104 59900 6 wbs_sel_i[1]
port 414 nsew signal input
rlabel metal2 s 43344 100 43400 400 6 wbs_sel_i[2]
port 415 nsew signal input
rlabel metal3 s 100 13104 400 13160 6 wbs_sel_i[3]
port 416 nsew signal input
rlabel metal3 s 100 49728 400 49784 6 wbs_stb_i
port 417 nsew signal input
rlabel metal3 s 59600 29232 59900 29288 6 wbs_we_i
port 418 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 11047988
string GDS_FILE /home/runner/work/RISCV-with-CNN-co-processor/RISCV-with-CNN-co-processor/openlane/tiny_user_project/runs/22_12_03_06_26/results/signoff/tiny_user_project.magic.gds
string GDS_START 345920
<< end >>

